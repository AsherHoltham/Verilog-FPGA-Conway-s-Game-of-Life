// global_variables.vh
