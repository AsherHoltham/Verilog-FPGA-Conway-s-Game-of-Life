`timescale 1ns / 1ps

module Game_of_Life;


endmodule