module set_up 
    (
        input integer death_cnt;
        input integer birth_cnt;
        input reg[0:0] input_board[15:0][15:0], 
        output reg[0:0] output_board[15:0][15:0]
    );


endmodule