module set_up 
    (
        input integer death_cnt;
        input integer birth_cnt;
        input environment_t input_environment, 
        output environment_t output_engironment
    );


endmodule