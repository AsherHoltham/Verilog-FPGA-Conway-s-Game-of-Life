// environment.vh
`ifndef ENVIRONMENT
`define ENVIRONMENT

// parameters
`define ENV_rows 16
`define ENV_cols 16

typedef bit [0:0] environment_t [`ENV_rows-1:0][`ENV_cols-1:0];

`endif