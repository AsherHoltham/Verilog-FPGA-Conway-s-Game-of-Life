// environment.vh
`ifndef ENVIRONMENT
`define ENVIRONMENT

typedef bit [0:0] environment_t [15:0][15:0];

`endif