module update_vga
    (

    );
    
endmodule