`timescale 1ns / 1ps

module vga_t
    (

    );

endmodule