module update_board_output 
    (

    );
    
endmodule